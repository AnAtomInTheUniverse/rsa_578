`ifdef DEFINES
`else
`define CLOCK_PERIOD 10  // DO NOT CHANGE
`define DEFINES 1
`define BITS 32
`define LOG_BITS 5
`endif
